`timescale 1ns/1ns

// ------------------------
// 6-by-6 unsigned fxp mult
// ------------------------

module mul_fp52 (
 clk
,op_a_dat	//|< r
,op_b_dat   //|< r
,op_c_dat   //|< r
,op_a_exp
,op_b_exp
,op_c_exp
,res
 );

input               clk;
input    [5:0] op_a_dat;  // 6-bit fraction: implicit + 5-bit mantissa + 1
input    [5:0] op_b_dat;
input    [5:0] op_c_dat;
input    [1:0] op_a_exp;  // 2-bit exponent
input    [1:0] op_b_exp;
input    [1:0] op_c_exp;
output  [17:0] res;       //12 + max(3+3,3) = 18 bits

reg    	 [5:0] op_a_dat_reg;
reg    	 [5:0] op_b_dat_reg;
reg    	 [5:0] op_c_dat_reg;
reg    	 [1:0] op_a_exp_reg;
reg    	 [1:0] op_b_exp_reg;
reg    	 [1:0] op_c_exp_reg;
wire   	[19:0] res_wire;
reg    	[19:0] res;

always@(posedge clk)
begin
    op_a_dat_reg <= op_a_dat;				
    op_b_dat_reg <= op_b_dat;
    op_c_dat_reg <= op_c_dat;
    op_a_exp_reg <= op_a_exp;				
    op_b_exp_reg <= op_b_exp;	
    op_c_exp_reg <= op_c_exp;	
    res 		 <= res_wire;
end

	mul u_mul( 
     .op_a_dat(op_a_dat_reg)
    ,.op_b_dat(op_b_dat_reg)
    ,.op_c_dat(op_c_dat_reg)
    ,.op_a_exp(op_a_exp_reg)
    ,.op_b_exp(op_b_exp_reg)
    ,.op_c_exp(op_c_exp_reg)
	,.res(res_wire)
    ,.clk(clk)
	);
endmodule   // wrapper

module mul (
 op_a_dat	//|< r
,op_b_dat	//|< r
,op_c_dat	//|< r
,op_a_exp
,op_b_exp
,op_c_exp
,res
,clk
 );

input               clk;
input    [5:0] op_a_dat;  // 6-bit fraction: implicit + 5-bit mantissa + 1
input    [5:0] op_b_dat;
input    [5:0] op_c_dat;
input    [1:0] op_a_exp;  // 2-bit exponent
input    [1:0] op_b_exp;
input    [1:0] op_c_exp;
output  [17:0] res;       //12 + max(3+3,3) = 18 bits

wire     [6:0] sel_data_0;
wire     [6:0] sel_data_1;
wire     [6:0] sel_data_2;
wire     [6:0] sel_data_3;
wire           sel_inv_0;
wire           sel_inv_1;
wire           sel_inv_2;
wire           sel_inv_3;

reg      [8:0] code_lo;
reg      [2:0] code_0;
reg      [2:0] code_1;
reg      [2:0] code_2;
reg      [2:0] code_3;

reg     [17:0] ppre_0;
reg     [17:0] ppre_1;
reg     [17:0] ppre_2;
reg     [17:0] ppre_3;
reg     [17:0] ppre_4;
reg     [17:0] ppre_5;

reg     [2:0] exp_sft;

reg     [17:0] ppre_0_sft;
reg     [17:0] ppre_1_sft;
reg     [17:0] ppre_2_sft;
reg     [17:0] ppre_3_sft;
reg     [17:0] ppre_4_sft;
reg     [17:0] ppre_5_sft;
reg     [17:0] ppre_6_sft;

reg     [53:0] pp_in_l0n0;
reg     [53:0] pp_in_l0n1;
wire    [17:0] pp_out_l0n0_0;
wire    [17:0] pp_out_l0n0_1;
wire    [17:0] pp_out_l0n1_0;
wire    [17:0] pp_out_l0n1_1;

reg     [89:0] pp_in_l1n0;
wire    [17:0] pp_out_l1n0_0;
wire    [17:0] pp_out_l1n0_1;

reg     [17:0] res;
//==========================================================
// Booth recoding and selection, radix-4
//==========================================================
always @(
	op_b_dat
  ) begin
    code_lo = {2'b0, op_b_dat, 1'b0};   // 9 bits
    code_0 = code_lo[2:0];
    code_1 = code_lo[4:2];
    code_2 = code_lo[6:4];
    code_3 = code_lo[8:6];
end

NV_NVDLA_CMAC_CORE_MAC_booth u_booth_0 (
   .code     (code_0[2:0])          //|< r
  ,.src_data (op_a_dat)   	        //|< r		
  ,.out_data (sel_data_0)           //|> w
  ,.out_inv  (sel_inv_0)            //|> w
  );

NV_NVDLA_CMAC_CORE_MAC_booth u_booth_1 (
   .code     (code_1[2:0])          //|< r
  ,.src_data (op_a_dat)  			//|< r
  ,.out_data (sel_data_1)           //|> w
  ,.out_inv  (sel_inv_1)            //|> w
  );
  
NV_NVDLA_CMAC_CORE_MAC_booth u_booth_2 (
   .code     (code_2[2:0])          //|< r
  ,.src_data (op_a_dat)   			//|< r
  ,.out_data (sel_data_2)           //|> w
  ,.out_inv  (sel_inv_2)            //|> w
  );

NV_NVDLA_CMAC_CORE_MAC_booth u_booth_3 (
   .code     (code_3[2:0])          //|< r
  ,.src_data (op_a_dat)   			//|< r
  ,.out_data (sel_data_3)           //|> w
  ,.out_inv  (sel_inv_3)            //|> w
  );

always @(
  sel_data_0
  or sel_data_1
  or sel_data_2
  or sel_data_3
  or sel_inv_0
  or sel_inv_1
  or sel_inv_2
  or sel_inv_3
  ) begin
    ppre_0 = {11'b0, sel_data_0};    // 18 bits
    ppre_1 = {9'b0, sel_data_1, 1'b0, sel_inv_0};
    ppre_2 = {7'b0, sel_data_2, 1'b0, sel_inv_1, 2'b0};
    ppre_3 = {5'b0, sel_data_3, 1'b0, sel_inv_2, 4'b0};
    ppre_4 = {11'b000_0000_0000, sel_inv_3, 6'b0};  // 1_1101_0101_1_000000
    ppre_5 = 18'b11_1110_1010_1100_0000;
end

always @(
    op_a_exp
    or op_b_exp
) begin
    exp_sft = op_a_exp + op_b_exp;
end

always @(
    ppre_0
    or ppre_1
    or ppre_2
) begin
    ppre_0_sft = ppre_0 << exp_sft;
    ppre_1_sft = ppre_1 << exp_sft;
    ppre_2_sft = ppre_2 << exp_sft;
end

always @(
    ppre_3
    or ppre_4
    or ppre_5
    or op_c_dat
    or op_c_exp
) begin
    ppre_3_sft = ppre_3 << exp_sft;
    ppre_4_sft = ppre_4 << exp_sft;
    ppre_5_sft = ppre_5 << exp_sft;
    ppre_6_sft = {12'b0, op_c_dat}<<op_c_exp;
end

//==========================================================
// CSA tree (level 1)
//==========================================================

always @(
    ppre_0_sft
    or ppre_1_sft
    or ppre_2_sft
    or ppre_3_sft
    or ppre_4_sft
    or ppre_5_sft
) begin
    pp_in_l0n0 = {ppre_2_sft, ppre_1_sft, ppre_0_sft};
    pp_in_l0n1 = {ppre_5_sft, ppre_4_sft, ppre_3_sft};
end

NV_DW02_tree #(3, 18) u_tree_l0n0 (							
   .INPUT    (pp_in_l0n0[53:0])      //|< r
  ,.OUT0     (pp_out_l0n0_0[17:0])   //|> sum
  ,.OUT1     (pp_out_l0n0_1[17:0])   //|> carry
  );
  
NV_DW02_tree #(3, 18) u_tree_l0n1 (							
   .INPUT    (pp_in_l0n1[53:0])      //|< r
  ,.OUT0     (pp_out_l0n1_0[17:0])   //|> sum
  ,.OUT1     (pp_out_l0n1_1[17:0])   //|> carry
  );

//==========================================================
// CSA tree (level 2)
//==========================================================
always @(
  /* pp_out_l0n1_1
  or pp_out_l0n1_0
  or pp_out_l0n0_1
  or pp_out_l0n0_0 */
  posedge clk
  ) begin
    pp_in_l1n0 = {ppre_6_sft, pp_out_l0n1_1, pp_out_l0n1_0, pp_out_l0n0_1, pp_out_l0n0_0};
end

NV_DW02_tree #(5, 18) u_tree_l1n0 (							
   .INPUT    (pp_in_l1n0[89:0])      //|< r
  ,.OUT0     (pp_out_l1n0_0[17:0])   //|> sum
  ,.OUT1     (pp_out_l1n0_1[17:0])   //|> carry
  );

always @(
    pp_out_l1n0_0
    or pp_out_l1n0_1
) begin
    res = pp_out_l1n0_1 + pp_out_l1n0_0;
end

endmodule // mul

//==========================================================
//
// Sub unit for mul
// Booth's recoder and Booth's selector with inversed sign flag
//
//==========================================================
module NV_NVDLA_CMAC_CORE_MAC_booth (
   code
  ,src_data
  ,out_data
  ,out_inv
  );

input    [2:0] code;
input    [5:0] src_data;
output   [6:0] out_data;
output         out_inv;

reg      [2:0] in_code;
reg      [6:0] out_data;
reg            out_inv;

always @(
  code
  or src_data
  ) begin
    case(code)
        ///////// for 6 bit /////////
        // +/- 0*src_data
        3'b000,
        3'b111:
        begin
            out_data = 7'b100_0000;
            out_inv = 1'b0;
        end

        // + 1*src_data
        3'b001,
        3'b010:
        begin
            out_data = {~src_data[5], src_data};
            out_inv = 1'b0;
        end

        // - 1*src_data
        3'b101,
        3'b110:
        begin
            out_data = {src_data[5], ~src_data};
            out_inv = 1'b1;
        end

        // + 2*src_data
        3'b011:
        begin
            out_data = {~src_data[5], src_data[4:0], 1'b0};	//shift
            out_inv = 1'b0;
        end

        // - 2*src_data
        3'b100:
        begin
            out_data = {src_data[5], ~src_data[4:0], 1'b1};	//shift and add
            out_inv = 1'b1;
        end
		
		default:
        begin
            out_data = 7'b100_0000;
            out_inv = 1'b0;
        end
    endcase
end
endmodule // NV_NVDLA_CMAC_CORE_MAC_booth